* RC_filter

*Sheet Name:/
R1  0 /n1 1k
C1  /n0 /n1 3.3nF		
V1  /n0 0 SIN(0 10 1kHz)		

.end
